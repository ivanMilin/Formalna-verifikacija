bind sv_model top c0(.clk(clk), .rst(rst), .x(x), .y(y));
