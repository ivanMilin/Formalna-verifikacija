bind and_case and_checker c0(.clk(clk), .rst(rst), .a(a), .b(b), .c(c));
bind and_wire and_checker c1(.clk(clk), .rst(rst), .a(a), .b(b), .c(c));
bind and_proc and_checker c2(.clk(clk), .rst(rst), .a(a), .b(b), .c(c));
